module CLK_Divider (input CLK,
						  output T_CLK);
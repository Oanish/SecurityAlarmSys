module Audio_Controller;

endmodule 
module Alarm_Controller(input CLK,					//trigger clock, used in all modules and by the DAC decoder
								input [7:0] Distance,	//distance from object, bits
								output Sound);				//alarm data stream to be converted to analog audio
								
//do stuff here

endmodule 
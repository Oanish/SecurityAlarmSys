module Sensor_Controller;

//IS NOT FINISHED